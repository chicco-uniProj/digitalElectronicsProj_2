library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



package costanti is
constant nbit: integer:=8;
end package costanti;